`include "definitions.v"
`timescale 1ns / 1ps

/*
this module handles hazards and interrupts 
 */

module hazard_unit (
    input clk, rst_n,

    input      uart_complete,                                   // from uart_unit (upg_done_i)
    output reg uart_disable,                                    // for (1) uart_unit (upg_rst_i)
                                                                //     (2) instruction_mem (switch to uart write mode)
                                                                //     (3) data_mem (switch to uart write mode)

    input      reg_1_valid,                                     // from signal_mux (whether register 1 is valid)
    input      reg_2_valid,                                     // from signal_mux (whether register 2 is valid)
    input      branch_instruction,                              // from control_unit (whether it is a branch instruction)

    input      ex_mem_read_enable,                              // from id_ex_reg (instruction needs to read from memory)
    input      ex_reg_write_enable,                             // from id_ex_reg (instruction needs write to register)
    input      ex_no_op,                                        // from id_ex_reg (the ex stage is a bubble)
    input      mem_reg_write_enable,                            // from ex_mem_reg (instruction needs write to register)
    input      mem_no_op,                                       // from ex_mem_reg (the mem stage is a bubble)

    input      [`REG_FILE_ADDR_WIDTH - 1:0] id_reg_1_idx,       // from signal_mux (index of first source register)
    input      [`REG_FILE_ADDR_WIDTH - 1:0] id_reg_2_idx,       // from signal_mux (index of second source register)
    input      [`REG_FILE_ADDR_WIDTH - 1:0] ex_reg_dest_idx,    // from id_ex_reg (index of destination resgiter)
    input      [`REG_FILE_ADDR_WIDTH - 1:0] mem_reg_dest_idx,   // from ex_mem_reg (index of destination resgiter)

    input      [`ISA_WIDTH - 1:0] pc_next,                      // from instruction_mem 

    input      input_enable,                                    // from data_mem (the keypad input is needed)
    input      input_complete,                                  // from keypad_unit (user pressed enter)
    input      cpu_pause,                                       // from keypad_unit (user pressed pause)

    output reg pc_reset,                                        // for instruction_mem (reset the pc to 0)
    output reg [1:0] if_hazard_control,                         // hazard control signal for each stage register
                     id_hazard_control,
                     ex_hazard_control,
                     mem_hazard_control,
                     wb_hazard_control,       
    output reg [2:0] issue_type                                 // for vga_unit (both hazard and interrupt)
    );
    
    reg [1:0] cpu_state;    // the state CPU is in

    wire mem_conflict = mem_reg_write_enable & ~mem_no_op &                     // wirte enabled and operational
                        ((reg_1_valid & id_reg_1_idx == mem_reg_dest_idx) |     // valid and conflict
                         (reg_2_valid & id_reg_2_idx == mem_reg_dest_idx));     // valid and conflict
    wire ex_conflict  = ex_reg_write_enable  & ~ex_no_op  &                     // wirte enabled and operational
                        ((reg_1_valid & id_reg_1_idx == ex_reg_dest_idx)  |     // valid and conflict
                         (reg_2_valid & id_reg_2_idx == ex_reg_dest_idx));      // valid and conflict
    
    wire data_hazard    = (branch_instruction & (ex_conflict | mem_conflict)) |     // data hazard when branch depends on data from previous stages 
                          (ex_mem_read_enable & ex_conflict);                       // data hazard when alu depends on data from memory at the next stage
    wire uart_hazard    = `PC_MAX_VALUE < pc_next;                                  // next instruction not in instruction memory

    wire data_resolved    = issue_type == `DATA   & ~data_hazard;
    wire uart_resolved    = issue_type == `UART   & uart_complete;
    wire pause_resolved   = issue_type == `PAUSE  & ~cpu_pause;

    always @(negedge clk, negedge rst_n) begin
        if (~rst_n) begin
            cpu_state    <= `IDLE;
            issue_type   <= `NONE;
            pc_reset     <= 1'b0;
            uart_disable <= 1'b1;
            {
                if_hazard_control, 
                id_hazard_control,
                ex_hazard_control,
                mem_hazard_control,
                wb_hazard_control
            }            <= 0;
        end else begin
            case (cpu_state) 
                `EXECUTE: begin
                    pc_reset     <= 1'b0;
                    casex ({data_hazard, cpu_pause, uart_hazard, input_enable})
                        // data hazard will hold all stages hence covers the other hazards
                        4'b1xxx: begin
                            issue_type <= `DATA;
                            // cpu_state  <= `HAZARD;
                            if_hazard_control <= `HOLD;  // if stage will not be a bubble
                            id_hazard_control <= `HOLD; // ex stage will be a bubble (the instruction in ex will enter wb by then)
                            ex_hazard_control <= `NO_OP;
                            // mem_hazard_control <= `;
                            // ex_hazard_control <= `NO_OP; // id stage will not be a bubble
                        end
                        // the user paused the CPU, the user can do UART rewrite during this period
                        4'b01xx: begin
                            issue_type   <= `PAUSE;
                            cpu_state    <= `HAZARD;
                            uart_disable <= 1'b0;
                            if_hazard_control <= `NO_OP; // start pumping no_op signals into the pipeline
                            id_hazard_control <= `NORMAL;
                        end
                        // the user did not pause the CPU but the pc overflowed, the CPU will automatically resume upon UART completion
                        4'b001x: begin
                            issue_type   <= `UART;
                            cpu_state    <= `HAZARD;
                            uart_disable <= 1'b0;
                            if_hazard_control <= `NO_OP;
                            id_hazard_control <= `NORMAL;
                        end
                        // CPU waits for the user's keypad input
                        4'b0001: begin
                            issue_type   <= `KEYPAD;
                            cpu_state    <= `INTERRUPT;
                            if_hazard_control   <= `NO_OP;
                            id_hazard_control   <= `NO_OP;
                            ex_hazard_control   <= `NO_OP;
                            mem_hazard_control  <= `NO_OP;
                            wb_hazard_control   <= `NO_OP;
                        end
                        default: begin
                            if_hazard_control   <= `NORMAL;
                            id_hazard_control   <= `NORMAL;
                            ex_hazard_control   <= `NORMAL;
                            mem_hazard_control  <= `NORMAL; 
                            wb_hazard_control   <= `NORMAL;
                        end
                    endcase
                end
                `HAZARD: begin
                    casex ({data_resolved, uart_resolved, pause_resolved})
                        3'b100 : begin
                            issue_type   <= `NONE;
                            cpu_state    <= `EXECUTE;
                            if_hazard_control   <= `NORMAL;
                            id_hazard_control   <= `NORMAL;
                            // ex_hazard_control   <= `NORMAL;
                        end
                        3'b01x : begin
                            issue_type   <= `PAUSE;
                            uart_disable <= 1'b1;
                            pc_reset     <= 1'b1;
                        end
                        3'b001 : begin
                            issue_type   <= `NONE;
                            cpu_state    <= `EXECUTE;
                            uart_disable <= 1'b1;
                            if_hazard_control   <= `NORMAL; // resuming the entire cpu from the next instruction
                        end
                        default: 
                            if (issue_type == `UART & (cpu_pause | uart_complete)) 
                                issue_type <= `PAUSE;       // pause after pc overflow which then the CPU must wait for the user to resume it
                            else 
                                issue_type <= issue_type;   // prevent auto latches
                    endcase
                end   
                `INTERRUPT: begin
                    if (input_complete) begin
                        issue_type <= `NONE;
                        cpu_state  <= `EXECUTE;
                        if_hazard_control   <= `RESUME;
                        id_hazard_control   <= `RESUME;
                        ex_hazard_control   <= `RESUME;
                        mem_hazard_control  <= `RESUME; 
                        wb_hazard_control   <= `RESUME;
                    end else 
                        issue_type <= issue_type; // prevent auto latches
                end
                default: // this is for `IDLE state, preventing auto latches
                    cpu_state <= `EXECUTE;
            endcase   
        end
    end
endmodule