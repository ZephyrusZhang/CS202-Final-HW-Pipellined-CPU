`timescale 1ns / 1ps

module seg_top ();



endmodule