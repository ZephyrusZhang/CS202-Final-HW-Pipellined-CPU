`timescale 1ns / 1ps

module top(
    input wire clk, rst_n,
    input wire [3:0] row_in,

    output reg [3:0] col_out
    output reg []

);
endmodule